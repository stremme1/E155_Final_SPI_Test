`timescale 1ns / 1ps

module spi_test_top (
    input  logic        fpga_rst_n,  // Global FPGA reset pin (active low)
    
    // SPI Interface (matches Sensor 1 in drum_set_top)
    output logic        sclk1,
    output logic        mosi1,
    input  logic        miso1,
    output logic        cs_n1,
    output logic        ps0_1,  // Added PS0/WAKE pin
    output logic        bno085_rst_n1, // BNO085 Reset pin (active low)
    input  logic        int1,
    
    // Button Inputs (EXACT from C code)
    input  logic        calibrate_btn_n,  // Button 2: Calibration (active low, with pull-up)
    input  logic        kick_btn_n,       // Button 1: Kick drum (active low, with pull-up)
    
    // Drum Trigger Outputs
    output logic        drum_trigger_valid,
    output logic [3:0]  drum_code,       // 0-7 (matches C code exactly)
    output logic        drum_hand,        // 0=right, 1=left
    
    // Debug / Status LEDs
    output logic        led_initialized, // ON when BNO085 init complete
    output logic        led_error,       // ON if error state
    output logic        led_heartbeat    // Blinks to show clock is running
);

    // Internal signals
    logic clk;
    logic rst_n;  // Internal reset signal
    logic spi_start, spi_tx_valid, spi_tx_ready, spi_rx_valid, spi_busy;
    logic [7:0] spi_tx_data, spi_rx_data;
    logic quat_valid, gyro_valid;
    logic signed [15:0] quat_w, quat_x, quat_y, quat_z;
    logic signed [15:0] gyro_x, gyro_y, gyro_z;
    logic initialized, error;
    
    // BNO085 Reset Delay Counter
    // Per datasheet 6.5.3: After NRST release, BNO085 needs:
    //   - t1 = 90ms for internal initialization
    //   - t2 = 4ms for internal configuration  
    //   - Total: ~94ms minimum, we use 100ms for safety
    // Clock is 3MHz, so 100ms = 300,000 cycles
    // We add 2 seconds total delay as requested
    localparam [22:0] DELAY_100MS = 23'd300_000;  // 100ms for BNO085 initialization
    localparam [22:0] DELAY_2SEC = 23'd6_000_000;  // 2 seconds total delay
    logic [22:0] rst_delay_counter;
    logic bno085_rst_n_delayed;
    logic controller_rst_n;  // Controller reset synchronized with BNO085 reset
    
    // BNO085 Reset with delay after FPGA reset release
    // Per datasheet 6.5.3: BNO085 needs ~94ms after NRST release before ready
    // Sequence: FPGA reset releases -> wait 100ms -> release BNO085 reset -> wait 1.9s -> release controller reset
    always_ff @(posedge clk or negedge fpga_rst_n) begin
        if (!fpga_rst_n) begin
            // FPGA reset is active: keep BNO085 in reset and reset counter
            rst_delay_counter <= 23'd0;
            bno085_rst_n_delayed <= 1'b0;
            controller_rst_n <= 1'b0;  // Keep controller in reset too
        end else begin
            // FPGA reset released: count up to delay
            if (rst_delay_counter < DELAY_2SEC) begin
                rst_delay_counter <= rst_delay_counter + 1;
            end
            
            // Release BNO085 reset after 100ms (allows BNO085 to initialize per datasheet)
            if (rst_delay_counter >= DELAY_100MS) begin
                bno085_rst_n_delayed <= 1'b1;  // Release BNO085 reset
            end else begin
                bno085_rst_n_delayed <= 1'b0;  // Keep BNO085 in reset
            end
            
            // Release controller reset after full 2-second delay
            // This ensures BNO085 has completed initialization before controller starts
            if (rst_delay_counter >= DELAY_2SEC) begin
                controller_rst_n <= 1'b1;  // Release controller reset
            end else begin
                controller_rst_n <= 1'b0;  // Keep controller in reset
            end
        end
    end
    
    assign bno085_rst_n1 = bno085_rst_n_delayed;
    assign rst_n = controller_rst_n;  // Controller reset synchronized with BNO085 reset release

    // HARDWARE CLOCK - HSOSC (ACTIVE FOR HARDWARE)
    // CLKHF_DIV(2'b11) = divide by 16 to get 3MHz from 48MHz
    // For 48MHz HSOSC: divide by 16 = 3MHz (suitable for SPI)
    // For different frequencies, adjust CLKHF_DIV:
    //   2'b00 = divide by 2
    //   2'b01 = divide by 4  
    //   2'b10 = divide by 8
    //   2'b11 = divide by 16
    
    // HARDWARE CLOCK - HSOSC (ACTIVE FOR HARDWARE)
    // Note: HSOSC is a built-in primitive for iCE40UP5k
    // Make sure your synthesis tool recognizes this primitive
    HSOSC #(.CLKHF_DIV(2'b11)) hf_osc (
        .CLKHFPU(1'b1),   // Power up (must be 1)
        .CLKHFEN(1'b1),   // Enable (must be 1)
        .CLKHF(clk)       // Output clock (3MHz from 48MHz / 16)
    );

    // Heartbeat LED (1Hz approx)
    // 3MHz = 3,000,000 cycles/sec. 2^22 = ~4M. Bit 21 toggles every ~0.7s
    logic [21:0] heartbeat_cnt;
    always_ff @(posedge clk or negedge rst_n) begin
        if (!rst_n) heartbeat_cnt <= 0;
        else heartbeat_cnt <= heartbeat_cnt + 1;
    end
    assign led_heartbeat = heartbeat_cnt[21];

    // SPI Master
    spi_master #(.CLK_DIV(2)) spi_master_inst (
        .clk(clk),
        .rst_n(rst_n),
        .start(spi_start),
        .tx_valid(spi_tx_valid),
        .tx_data(spi_tx_data),
        .tx_ready(spi_tx_ready),
        .rx_valid(spi_rx_valid),
        .rx_data(spi_rx_data),
        .busy(spi_busy),
        .sclk(sclk1),
        .mosi(mosi1),
        .miso(miso1)
    );

    // BNO085 Controller
    bno085_controller bno085_ctrl_inst (
        .clk(clk),
        .rst_n(rst_n),
        .spi_start(spi_start),
        .spi_tx_valid(spi_tx_valid),
        .spi_tx_data(spi_tx_data),
        .spi_tx_ready(spi_tx_ready),
        .spi_rx_valid(spi_rx_valid),
        .spi_rx_data(spi_rx_data),
        .spi_busy(spi_busy),
        .cs_n(cs_n1),
        .ps0_wake(ps0_1),
        .int_n(int1),
        .quat_valid(quat_valid),
        .quat_w(quat_w),
        .quat_x(quat_x),
        .quat_y(quat_y),
        .quat_z(quat_z),
        .gyro_valid(gyro_valid),
        .gyro_x(gyro_x),
        .gyro_y(gyro_y),
        .gyro_z(gyro_z),
        .initialized(initialized),
        .error(error)
    );

    // Status LEDs
    assign led_initialized = initialized;
    assign led_error = error;
    
    // Button Debouncers (EXACT from C code: 50ms debounce)
    logic calibrate_btn_pulse, kick_btn_pulse;
    
    button_debouncer #(.DEBOUNCE_CYCLES(150000)) calibrate_debouncer (
        .clk(clk),
        .rst_n(rst_n),
        .btn_n(calibrate_btn_n),
        .btn_pressed(calibrate_btn_pulse),
        .btn_released(),
        .btn_state()
    );
    
    button_debouncer #(.DEBOUNCE_CYCLES(150000)) kick_debouncer (
        .clk(clk),
        .rst_n(rst_n),
        .btn_n(kick_btn_n),
        .btn_pressed(kick_btn_pulse),
        .btn_released(),
        .btn_state()
    );
    
    // Drum Trigger Processor
    drum_trigger_processor drum_processor (
        .clk(clk),
        .rst_n(rst_n),
        .quat1_valid(quat_valid),
        .quat1_w(quat_w),
        .quat1_x(quat_x),
        .quat1_y(quat_y),
        .quat1_z(quat_z),
        .gyro1_valid(gyro_valid),
        .gyro1_x(gyro_x),
        .gyro1_y(gyro_y),
        .gyro1_z(gyro_z),
        .calibrate_btn_pulse(calibrate_btn_pulse),
        .kick_btn_pulse(kick_btn_pulse),
        .drum_trigger_valid(drum_trigger_valid),
        .drum_code(drum_code),
        .drum_hand(drum_hand)
    );

endmodule
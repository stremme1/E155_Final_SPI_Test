Warning	1026001	Project	WARNING <1026001> - C:/Users/estralka/Desktop/E155_11.26/Final_FPGA_11_26/Ass_1.pdc (1) : No port matched 'miso_mcu'. [Ass_1.pdc:1]	
Warning	35935050	Synthesis	WARNING <35935050> - input port TRIM9 is not connected on this instance. VDB-5050	
Info	35901328	Synthesis	INFO <35901328> - c:/lscc/radiant/2024.2/ip/pmi/pmi_ice40up.v(1): analyzing included file c:/lscc/radiant/2024.2/ip/pmi/pmi_addsub.v. VERI-1328 [pmi_ice40up.v:1]	
Info	35921014	Synthesis	INFO <35921014> - c:/lscc/radiant/2024.2/ip/pmi/pmi_ice40up.vhd(4): analyzing package components. VHDL-1014 [pmi_ice40up.vhd:4]	
Info	35921504	Synthesis	INFO <35921504> - The default VHDL library search path is now "C:/Users/estralka/Desktop/E155_11.26/Final_FPGA_11_26/impl_1". VHDL-1504	
Info	35901018	Synthesis	INFO <35901018> - c:/users/estralka/desktop/e155_11.26/fpga/drum_trigger_top.sv(15): compiling module drum_trigger_top. VERI-1018 [drum_trigger_top.sv:15]	
Warning	35901209	Synthesis	WARNING <35901209> - c:/users/estralka/desktop/e155_11.26/fpga/drum_trigger_top.sv(83): expression size 32 truncated to fit in target size 23. VERI-1209 [drum_trigger_top.sv:83]	
Warning	35935040	Synthesis	WARNING <35935040> - Register \spi_slave_mcu_inst/shift_started_2 clock is stuck at Zero. VDB-5040	
Info	35001774	Synthesis	INFO <35001774> - Extracted state machine for register '\spi_master_inst1/state' with one-hot encoding	
Warning	35001714	Synthesis	WARNING <35001714> - Net gnd has following drivers :	
Error	35931000	Synthesis	ERROR <35931000> - c:/users/estralka/desktop/e155_11.26/fpga/spi_slave_mcu.sv(135): net gnd is constantly driven from multiple places at instance \spi_slave_mcu_inst/shift_started, on port q. VDB-1000 [spi_slave_mcu.sv:135]	
Project (16 warnings)	
Synthesis (1 errors, 4 criticals, 28 warnings, 41 info)	



`timescale 1ns / 1ps

// MCU SPI Slave Module
// FPGA is SPI slave to MCU (MCU is master) - READ-ONLY MODE
// Sends RAW sensor data packets to MCU
// Based on e155-lab7-main 2/fpga/src/aes_spi.sv pattern
// SPI Mode 0 (CPOL=0, CPHA=0): MCU samples on rising edge, FPGA changes on falling edge
// 
// Read-Only Protocol:
// - FPGA ignores MOSI (sdi) completely - only shifts out data on MISO (sdo)
// - MCU generates SCK by sending dummy bytes (0x00) via spiSendReceive(0)
// - FPGA shifts out 1 bit per SCK edge from its shift register
// - MCU reads data from MISO during the transaction

module spi_slave_mcu(
    input  logic        clk,           // FPGA system clock
    input  logic        sck,           // SPI clock from MCU (generated by MCU)
    input  logic        sdi,           // SPI data in (MOSI from MCU - IGNORED in read-only mode)
    output logic        sdo,           // SPI data out (MISO to MCU - shifts out data)
    input  logic        cs_n,          // Chip select from MCU (active low: CS low = transaction active)
    input  logic        load,          // Load signal from MCU (not used in simple CS pattern)
    output logic        done,          // Done signal to MCU (not used in simple CS pattern)
    
    // Sensor data inputs (RAW data from BNO085 controller)
    // Sensor 1 (Right Hand) - Single sensor only
    input  logic        quat1_valid,
    input  logic signed [15:0] quat1_w, quat1_x, quat1_y, quat1_z,
    input  logic        gyro1_valid,
    input  logic signed [15:0] gyro1_x, gyro1_y, gyro1_z
);

    // Packet format: 16 bytes total (single sensor only)
    // Byte 0:    Header (0xAA)
    // Byte 1-8:  Sensor 1 Quaternion (w, x, y, z - MSB,LSB each)
    // Byte 9-14: Sensor 1 Gyroscope (x, y, z - MSB,LSB each)
    // Byte 15:   Sensor 1 Flags (bit 0=quat_valid, bit 1=gyro_valid)
    
    localparam PACKET_SIZE = 16;
    localparam HEADER_BYTE = 8'hAA;
    
    // Packet buffer - assembled from sensor data
    logic [7:0] packet_buffer [0:PACKET_SIZE-1];
    logic       sdodelayed;  // Delayed SDO output for SPI Mode 0 timing
    
    // Assemble packet from sensor data (using assign statements for iverilog compatibility)
    // Header
    assign packet_buffer[0] = HEADER_BYTE;
    
    // Sensor 1 Quaternion (MSB,LSB format)
    assign packet_buffer[1] = quat1_w[15:8];  // W MSB
    assign packet_buffer[2] = quat1_w[7:0];   // W LSB
    assign packet_buffer[3] = quat1_x[15:8];  // X MSB
    assign packet_buffer[4] = quat1_x[7:0];   // X LSB
    assign packet_buffer[5] = quat1_y[15:8];  // Y MSB
    assign packet_buffer[6] = quat1_y[7:0];   // Y LSB
    assign packet_buffer[7] = quat1_z[15:8];  // Z MSB
    assign packet_buffer[8] = quat1_z[7:0];   // Z LSB
    
    // Sensor 1 Gyroscope (MSB,LSB format)
    assign packet_buffer[9]  = gyro1_x[15:8];  // X MSB
    assign packet_buffer[10] = gyro1_x[7:0];   // X LSB
    assign packet_buffer[11] = gyro1_y[15:8];  // Y MSB
    assign packet_buffer[12] = gyro1_y[7:0];   // Y LSB
    assign packet_buffer[13] = gyro1_z[15:8];  // Z MSB
    assign packet_buffer[14] = gyro1_z[7:0];   // Z LSB
    
    // Sensor 1 Flags
    assign packet_buffer[15] = {6'h0, gyro1_valid, quat1_valid};
    
    // Simple CS-based pattern: Use CS to detect transaction boundaries
    // FPGA always has latest packet_buffer data ready
    // Shift register is loaded when CS goes low (transaction starts)
    // DONE/LOAD signals not used in simple CS pattern
    assign done = 1'b1;  // Always ready - MCU doesn't check this in simple pattern
    
    // Create a 128-bit shift register from packet buffer (16 bytes * 8 bits)
    // Read-only mode: FPGA ignores MOSI (sdi), only shifts out data on MISO (sdo)
    // Simple CS-based pattern: Load on first SCK edge when CS is low, shift on subsequent SCK edges
    logic [127:0] packet_shift_reg;
    logic cs_n_prev_sck = 1'b1;  // Track previous CS state in SCK domain to detect falling edge
    
    // SPI Mode 0 (CPOL=0, CPHA=0): MCU samples on rising edge, FPGA changes on falling edge
    // Shift register behavior:
    // - On first posedge when CS is low: load latest packet_buffer into shift register
    // - On subsequent posedges when CS is low: shift left (MSB first) - FPGA ignores SDI (MOSI)
    // - All updates happen in SCK clock domain to avoid multiple drivers
    always_ff @(posedge sck) begin
        cs_n_prev_sck <= cs_n;  // Track CS state in SCK domain
        
        if (!cs_n) begin
            if (cs_n_prev_sck) begin
                // First SCK edge after CS went low: load latest packet buffer into shift register (MSB first)
                // Pack all bytes: packet_buffer[0] is MSB of first byte, goes to bit 127
                // Read-only mode: ignore SDI (MOSI), only shift out data
                // Always load latest data - no need to wait for done signal
                packet_shift_reg <= {
                    packet_buffer[0], packet_buffer[1], packet_buffer[2], packet_buffer[3],
                    packet_buffer[4], packet_buffer[5], packet_buffer[6], packet_buffer[7],
                    packet_buffer[8], packet_buffer[9], packet_buffer[10], packet_buffer[11],
                    packet_buffer[12], packet_buffer[13], packet_buffer[14], packet_buffer[15]
                };
            end else begin
                // Subsequent SCK edges: shift left (MSB first)
                // Read-only mode: ignore SDI, shift in 0 (or just shift left)
                packet_shift_reg <= {packet_shift_reg[126:0], 1'b0};
            end
        end
    end
    
    // Update output on negedge (when FPGA should change MISO for next bit)
    // Only update when CS is low (transaction active)
    always_ff @(negedge sck) begin
        if (!cs_n) begin
            // After shift on posedge, the new MSB is at bit 126 (bit 127 was shifted out)
            // This is the bit that will be sampled on the next posedge
            sdodelayed = packet_shift_reg[126];  // New MSB after shift
        end
    end
    
    // Track if we've started shifting (after first SCK edge)
    logic shift_started = 1'b0;
    
    // Reset shift_started when CS goes high (transaction ends)
    always_ff @(posedge clk) begin
        if (cs_n) begin
            shift_started <= 1'b0;  // CS is high, reset for next transaction
        end
    end
    
    // Set shift_started after first SCK edge
    always_ff @(posedge sck) begin
        if (!cs_n) begin
            shift_started <= 1'b1;  // First SCK edge in transaction
        end
    end
    
    // SDO (MISO) output: Read-only mode
    // SPI Mode 0 timing:
    // - When CS is high: output 0 (not in transaction)
    // - When CS is low and before first SCK edge: output MSB directly from packet_buffer[0][7]
    // - After first SCK edge: use sdodelayed (set on negedge)
    // packet_buffer[0][7] is MSB of first byte (bit 7 of byte 0), which is MSB of entire packet
    // sdodelayed is updated on negedge to packet_shift_reg[127] (current MSB)
    assign sdo = (!cs_n && !shift_started) ? packet_buffer[0][7] : 
                 (!cs_n) ? sdodelayed : 1'b0;  // Output 0 when CS is high (not selected)
    
endmodule



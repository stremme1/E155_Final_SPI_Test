`timescale 1ns / 1ps

// Comprehensive Testbench for BNO085 SPI Controller
// Tests:
// 1. PS0/WAKE sequence per datasheet
// 2. Initialization commands (Product ID, Rotation Vector, Gyroscope)
// 3. SHTP protocol compliance
// 4. Data report reading

module tb_spi_test;

    // Signal declarations matching spi_test_top
    logic rst_n;
    logic sclk1;
    logic mosi1;
    logic miso1;
    logic cs_n1;
    logic ps0_1;  // PS0/WAKE pin
    logic int1;
    logic led_initialized;
    logic led_error;
    logic led_heartbeat;

    // Instantiate the DUT (Device Under Test)
    spi_test_top dut (
        .rst_n(rst_n),
        .sclk1(sclk1),
        .mosi1(mosi1),
        .miso1(miso1),
        .cs_n1(cs_n1),
        .ps0_1(ps0_1),
        .int1(int1),
        .led_initialized(led_initialized),
        .led_error(led_error),
        .led_heartbeat(led_heartbeat)
    );

    // Instantiate the Mock BNO085 Sensor
    mock_bno085 sensor_model (
        .clk(dut.clk),
        .rst_n(rst_n),
        .ps0_wake(ps0_1),
        .cs_n(cs_n1),
        .sclk(sclk1),
        .mosi(mosi1),
        .miso(miso1),
        .int_n(int1)
    );

    // Test state tracking
    integer test_step = 0;
    integer init_commands_received = 0;
    logic [7:0] last_cmd_channel = 0;
    logic [7:0] last_cmd_seq = 0;

    // Accelerator: Skip long delays for faster simulation
    initial begin
        wait(rst_n == 1);
        forever begin
            @(posedge dut.clk);
            // INIT_WAIT_RESET: Skip most of 300,000 count delay
            if (dut.bno085_ctrl_inst.state == 1) begin // INIT_WAIT_RESET
                if (dut.bno085_ctrl_inst.delay_counter < 19'd299_900) begin
                    force dut.bno085_ctrl_inst.delay_counter = 19'd299_990;
                    @(posedge dut.clk);
                    release dut.bno085_ctrl_inst.delay_counter;
                end
            end
            // INIT_DONE_CHECK: Skip most of 30,000 count delay
            else if (dut.bno085_ctrl_inst.state == 5) begin // INIT_DONE_CHECK
                if (dut.bno085_ctrl_inst.delay_counter < 19'd29_900) begin
                    force dut.bno085_ctrl_inst.delay_counter = 19'd29_990;
                    @(posedge dut.clk);
                    release dut.bno085_ctrl_inst.delay_counter;
                end
            end
        end
    end

    // Monitor SPI transactions
    initial begin
        forever begin
            @(posedge cs_n1); // Wait for CS to go high (transaction end)
            #100;
            if (dut.bno085_ctrl_inst.state == 5) begin // INIT_DONE_CHECK
                init_commands_received = init_commands_received + 1;
                $display("[%0t] Command %0d completed", $time, init_commands_received);
            end
        end
    end

    // Main Test Sequence
    initial begin
        $dumpfile("spi_test.vcd");
        $dumpvars(0, tb_spi_test);

        $display("========================================");
        $display("BNO085 SPI Controller Testbench");
        $display("========================================");
        
        // 1. Reset System
        $display("\n[TEST] Step 1: System Reset");
        rst_n = 0;
        #1000;
        rst_n = 1;
        $display("[TEST] Reset released at %0t", $time);
        
        // Verify PS0 is high after reset (SPI mode selection)
        #100;
        if (ps0_1 == 1'b1) begin
            $display("[PASS] PS0 is HIGH after reset (SPI mode)");
        end else begin
            $display("[FAIL] PS0 should be HIGH after reset");
        end

        // 2. Wait for Initialization Sequence
        $display("\n[TEST] Step 2: Waiting for Initialization Sequence");
        $display("  - Product ID Request");
        $display("  - Enable Rotation Vector");
        $display("  - Enable Gyroscope");
        
        fork
            begin
                // Wait for initialized signal
                wait(dut.bno085_ctrl_inst.initialized == 1);
                $display("\n[PASS] Controller Initialized!");
                $display("  - LED status: %b", led_initialized);
                $display("  - Commands sent: %0d", init_commands_received);
                
                if (init_commands_received >= 3) begin
                    $display("[PASS] All 3 initialization commands completed");
                end else begin
                    $display("[FAIL] Expected 3 commands, got %0d", init_commands_received);
                end
            end
            begin
                // Timeout after 50ms simulation time
                #50000000; 
                $display("\n[FAIL] TIMEOUT waiting for initialization!");
                $display("  Current State: %0d", dut.bno085_ctrl_inst.state);
                $display("  Byte Count: %0d", dut.bno085_ctrl_inst.byte_cnt);
                $display("  INT_N: %b", int1);
                $display("  CS_N: %b", cs_n1);
                $display("  PS0: %b", ps0_1);
                $display("  Delay Counter: %0d", dut.bno085_ctrl_inst.delay_counter);
                $display("  CMD Select: %0d", dut.bno085_ctrl_inst.cmd_select);
                $finish;
            end
        join_any

        // 3. Test PS0 Wake Sequence
        $display("\n[TEST] Step 3: Verify PS0 Wake Sequence");
        // Controller should have used PS0 during init, verify it's released now
        if (ps0_1 == 1'b1) begin
            $display("[PASS] PS0 released after initialization");
        end else begin
            $display("[FAIL] PS0 should be HIGH in normal operation");
        end

        // 4. Test Rotation Vector Report
        $display("\n[TEST] Step 4: Testing Rotation Vector Report");
        #5000;
        
        // Send a test quaternion: W=1.0 (0x4000), X=0, Y=0, Z=0
        $display("  Sending Rotation Vector: W=0x4000, X=0, Y=0, Z=0");
        sensor_model.send_rotation_vector(16'd0, 16'd0, 16'd0, 16'h4000);
        
        fork
            begin
                wait(dut.bno085_ctrl_inst.quat_valid == 1);
                $display("\n[PASS] Quaternion Received!");
                $display("  W=%04h X=%04h Y=%04h Z=%04h", 
                         dut.bno085_ctrl_inst.quat_w, 
                         dut.bno085_ctrl_inst.quat_x, 
                         dut.bno085_ctrl_inst.quat_y, 
                         dut.bno085_ctrl_inst.quat_z);

                if (dut.bno085_ctrl_inst.quat_w == 16'h4000 &&
                    dut.bno085_ctrl_inst.quat_x == 16'd0 &&
                    dut.bno085_ctrl_inst.quat_y == 16'd0 &&
                    dut.bno085_ctrl_inst.quat_z == 16'd0) begin
                    $display("[PASS] Quaternion data matches expected values");
                end else begin
                    $display("[FAIL] Quaternion data mismatch");
                end
            end
            begin
                #2000000; // 2ms timeout
                $display("\n[FAIL] TIMEOUT waiting for quaternion data!");
                $finish;
            end
        join_any

        // 5. Test Gyroscope Report
        $display("\n[TEST] Step 5: Testing Gyroscope Report");
        #10000;
        
        // Send test gyro data: X=100, Y=200, Z=300
        $display("  Sending Gyroscope: X=100, Y=200, Z=300");
        sensor_model.send_gyroscope(16'd100, 16'd200, 16'd300);
        
        fork
            begin
                wait(dut.bno085_ctrl_inst.gyro_valid == 1);
                $display("\n[PASS] Gyroscope Received!");
                $display("  X=%04h Y=%04h Z=%04h", 
                         dut.bno085_ctrl_inst.gyro_x, 
                         dut.bno085_ctrl_inst.gyro_y, 
                         dut.bno085_ctrl_inst.gyro_z);

                if (dut.bno085_ctrl_inst.gyro_x == 16'd100 &&
                    dut.bno085_ctrl_inst.gyro_y == 16'd200 &&
                    dut.bno085_ctrl_inst.gyro_z == 16'd300) begin
                    $display("[PASS] Gyroscope data matches expected values");
                end else begin
                    $display("[FAIL] Gyroscope data mismatch");
                end
            end
            begin
                #2000000; // 2ms timeout
                $display("\n[FAIL] TIMEOUT waiting for gyroscope data!");
                $finish;
            end
        join_any

        // 6. Final Status Check
        $display("\n[TEST] Step 6: Final Status Check");
        if (led_error == 1'b0) begin
            $display("[PASS] Error LED is OFF");
        end else begin
            $display("[FAIL] Error LED is ON");
        end
        
        if (led_initialized == 1'b1) begin
            $display("[PASS] Initialized LED is ON");
        end else begin
            $display("[FAIL] Initialized LED is OFF");
        end

        #10000;
        $display("\n========================================");
        $display("All Tests Completed Successfully!");
        $display("========================================");
        $finish;
    end

    // Monitor for errors
    always @(posedge dut.bno085_ctrl_inst.error) begin
        $display("\n[ERROR] Controller entered error state at %0t", $time);
        $display("  State: %0d", dut.bno085_ctrl_inst.state);
    end

endmodule

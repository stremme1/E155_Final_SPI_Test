`timescale 1ns / 1ps

// MCU SPI Slave Module
// FPGA is SPI slave to MCU (MCU is master) - READ-ONLY MODE
// Sends RAW sensor data packets to MCU
// Based on e155-lab7-main 2/fpga/src/aes_spi.sv pattern
// SPI Mode 0 (CPOL=0, CPHA=0): MCU samples on rising edge, FPGA changes on falling edge
// 
// Read-Only Protocol:
// - FPGA ignores MOSI (sdi) completely - only shifts out data on MISO (sdo)
// - MCU generates SCK by sending dummy bytes (0x00) via spiSendReceive(0)
// - FPGA shifts out 1 bit per SCK edge from its shift register
// - MCU reads data from MISO during the transaction

module spi_slave_mcu(
    input  logic        clk,           // FPGA system clock
    input  logic        sck,           // SPI clock from MCU (generated by MCU)
    input  logic        sdi,           // SPI data in (MOSI from MCU - IGNORED in read-only mode)
    output logic        sdo,           // SPI data out (MISO to MCU - shifts out data)
    // Note: LOAD/DONE ports removed for CS-only operation
    
    // Sensor data inputs (RAW data from BNO085 controller)
    // Sensor 1 (Right Hand) - Single sensor only
    input  logic        quat1_valid,
    input  logic signed [15:0] quat1_w, quat1_x, quat1_y, quat1_z,
    input  logic        gyro1_valid,
    input  logic signed [15:0] gyro1_x, gyro1_y, gyro1_z
);

    // Packet format: 16 bytes total (single sensor only)
    // Byte 0:    Header (0xAA)
    // Byte 1-8:  Sensor 1 Quaternion (w, x, y, z - MSB,LSB each)
    // Byte 9-14: Sensor 1 Gyroscope (x, y, z - MSB,LSB each)
    // Byte 15:   Sensor 1 Flags (bit 0=quat_valid, bit 1=gyro_valid)
    
    localparam PACKET_SIZE = 16;
    localparam HEADER_BYTE = 8'hAA;
    
    // Packet buffer - assembled from sensor data
    logic [7:0] packet_buffer [0:PACKET_SIZE-1];
    logic       sdodelayed;
    logic       shift_reg_loaded = 1'b0;  // Track if shift register has been loaded in current transaction
    
    // Assemble packet from sensor data (using assign statements for iverilog compatibility)
    // Header
    assign packet_buffer[0] = HEADER_BYTE;
    
    // Sensor 1 Quaternion (MSB,LSB format)
    assign packet_buffer[1] = quat1_w[15:8];  // W MSB
    assign packet_buffer[2] = quat1_w[7:0];   // W LSB
    assign packet_buffer[3] = quat1_x[15:8];  // X MSB
    assign packet_buffer[4] = quat1_x[7:0];   // X LSB
    assign packet_buffer[5] = quat1_y[15:8];  // Y MSB
    assign packet_buffer[6] = quat1_y[7:0];   // Y LSB
    assign packet_buffer[7] = quat1_z[15:8];  // Z MSB
    assign packet_buffer[8] = quat1_z[7:0];   // Z LSB
    
    // Sensor 1 Gyroscope (MSB,LSB format)
    assign packet_buffer[9]  = gyro1_x[15:8];  // X MSB
    assign packet_buffer[10] = gyro1_x[7:0];   // X LSB
    assign packet_buffer[11] = gyro1_y[15:8];  // Y MSB
    assign packet_buffer[12] = gyro1_y[7:0];   // Y LSB
    assign packet_buffer[13] = gyro1_z[15:8];  // Z MSB
    assign packet_buffer[14] = gyro1_z[7:0];   // Z LSB
    
    // Sensor 1 Flags
    assign packet_buffer[15] = {6'h0, gyro1_valid, quat1_valid};
    
    // CS-only operation: Data is always available when valid sensor data is present
    // No LOAD/DONE handshaking needed - shift register loads on first SCK edge after idle
    
    // Create a 128-bit shift register from packet buffer (16 bytes * 8 bits)
    // Read-only mode: FPGA ignores MOSI (sdi), only shifts out data on MISO (sdo)
    logic [127:0] packet_shift_reg;
    
    // SPI Mode 0 (CPOL=0, CPHA=0): MCU samples on rising edge, FPGA changes on falling edge
    // CS-only operation: Shift register loads on first posedge, shifts on subsequent edges
    // Reset shift_reg_loaded when SCK has been idle (CS high) - detected on system clock
    always_ff @(posedge sck) begin
        if (!shift_reg_loaded) begin
            // First posedge after idle: load packet buffer into shift register (MSB first)
            // Pack all bytes: packet_buffer[0] is MSB of first byte, goes to bit 127
            // Read-only mode: ignore SDI (MOSI), only shift out data
            packet_shift_reg = {
                packet_buffer[0], packet_buffer[1], packet_buffer[2], packet_buffer[3],
                packet_buffer[4], packet_buffer[5], packet_buffer[6], packet_buffer[7],
                packet_buffer[8], packet_buffer[9], packet_buffer[10], packet_buffer[11],
                packet_buffer[12], packet_buffer[13], packet_buffer[14], packet_buffer[15]
            };
            shift_reg_loaded <= 1'b1;
        end else begin
            // Subsequent posedges: shift left (MSB first)
            // Read-only mode: ignore SDI, shift in 0
            packet_shift_reg = {packet_shift_reg[126:0], 1'b0};
        end
    end
    
    // Reset shift_reg_loaded when SCK has been idle (CS high)
    // Detect SCK idle by monitoring on system clock - if SCK stays low for many cycles, transaction is over
    logic sck_sync, sck_sync_prev;
    logic [7:0] sck_idle_counter = 8'd0;
    always_ff @(posedge clk) begin
        sck_sync <= sck;  // Synchronize SCK to system clock
        sck_sync_prev <= sck_sync;
        
        if (sck_sync && !sck_sync_prev) begin
            // SCK rising edge detected - reset idle counter
            sck_idle_counter <= 8'd0;
        end else if (!sck_sync) begin
            // SCK is low/idle - count up
            if (sck_idle_counter < 8'd255) begin
                sck_idle_counter <= sck_idle_counter + 1;
            end
            // If SCK has been idle for many cycles (>100), reset shift_reg_loaded for next transaction
            if (sck_idle_counter > 8'd100) begin
                shift_reg_loaded <= 1'b0;
            end
        end
    end
    
    // Update output on negedge (when FPGA should change MISO for next bit)
    // SPI Mode 0: FPGA changes MISO on falling edge, MCU samples on rising edge
    always_ff @(negedge sck) begin
        // After shift on posedge, next bit to output is at bit 126 (was at 127 before shift)
        sdodelayed = packet_shift_reg[126];  // Next bit to output (MSB of remaining data)
    end
    
    // SDO (MISO) output: Read-only mode, CS-only operation
    // SPI Mode 0 timing:
    // - Before first posedge: output MSB directly from packet_buffer[0][7]
    // - After first negedge: use sdodelayed (set on negedge)
    // packet_buffer[0][7] is MSB of first byte (bit 7 of byte 0), which is MSB of entire packet
    assign sdo = (!shift_reg_loaded) ? packet_buffer[0][7] : sdodelayed;
    
endmodule



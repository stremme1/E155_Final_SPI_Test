`timescale 1ns / 1ps

// Comprehensive Testbench for MCU SPI Slave Module (CS-based protocol)
// Tests SPI Mode 0 operation with CS control
// Verifies shift register behavior and packet transmission

module tb_spi_slave_mcu_debug;

    // Clock
    logic clk;
    
    // SPI interface (MCU is master, CS-based protocol)
    logic cs_n;      // Chip select from MCU (active low)
    logic sck;       // SPI clock from MCU
    logic sdi;       // SPI data in (MOSI - not used in read-only mode)
    logic sdo;       // SPI data out (MISO to MCU)
    
    // Sensor data inputs (single sensor only)
    logic quat1_valid, gyro1_valid;
    logic signed [15:0] quat1_w, quat1_x, quat1_y, quat1_z;
    logic signed [15:0] gyro1_x, gyro1_y, gyro1_z;
    
    // Clock generation (3MHz FPGA clock)
    parameter CLK_PERIOD = 333;
    always begin
        clk = 0;
        #(CLK_PERIOD/2);
        clk = 1;
        #(CLK_PERIOD/2);
    end
    
    // MCU SPI clock - NOT continuous! Only toggles during spiSendReceive calls
    // In real MCU, SCK only toggles when spiSendReceive() is called
    // SCK starts idle low (SPI Mode 0: CPOL=0)
    parameter SCK_PERIOD = 1000;  // 1MHz (1000ns period)
    initial begin
        sck = 0;  // Idle low for SPI Mode 0
    end
    // No continuous clock - SCK is controlled manually in tests
    
    // DUT
    spi_slave_mcu dut (
        .clk(clk),
        .cs_n(cs_n),
        .sck(sck),
        .sdi(sdi),
        .sdo(sdo),
        .initialized(1'b1),
        .error(1'b0),
        .quat1_valid(quat1_valid),
        .quat1_w(quat1_w),
        .quat1_x(quat1_x),
        .quat1_y(quat1_y),
        .quat1_z(quat1_z),
        .gyro1_valid(gyro1_valid),
        .gyro1_x(gyro1_x),
        .gyro1_y(gyro1_y),
        .gyro1_z(gyro1_z)
    );
    
    // Access internal signals for debugging
    wire [7:0] shift_out = dut.shift_out;
    wire [3:0] byte_count = dut.byte_count;
    wire [2:0] bit_count = dut.bit_count;
    wire [127:0] tx_packet = dut.tx_packet;
    
    // Access clock domain crossing and snapshot signals for debugging
    wire quat1_valid_snap = dut.quat1_valid_snap;
    wire gyro1_valid_snap = dut.gyro1_valid_snap;
    wire signed [15:0] quat1_w_snap = dut.quat1_w_snap;
    wire signed [15:0] quat1_x_snap = dut.quat1_x_snap;
    wire signed [15:0] gyro1_x_snap = dut.gyro1_x_snap;
    
    // Test variables
    logic [7:0] received_packet [0:15];
    integer test_count = 0;
    integer pass_count = 0;
    integer fail_count = 0;
    
    // Test loop variables
    integer bit_idx;
    logic sampled_bit;
    logic expected_bit;
    integer i, j;
    
    // Helper task to check and report
    task check_test(input string test_name, input logic condition);
        test_count = test_count + 1;
        if (condition) begin
            $display("[PASS] %s", test_name);
            pass_count = pass_count + 1;
        end else begin
            $display("[FAIL] %s", test_name);
            fail_count = fail_count + 1;
        end
    endtask
    
    // Task: MCU reads 16-byte packet via SPI Mode 0
    // SPI Mode 0: CPOL=0 (idle low), CPHA=0 (sample on rising edge)
    // Updated to properly simulate MCU SPI clock timing
    task mcu_read_packet_cs;
        integer i, j;
        logic [15:0] data_before_transaction;
        begin
            $display("[%0t] MCU: Starting SPI transaction - CS goes low", $time);
            
            // Capture data before transaction starts (for stability check)
            data_before_transaction = quat1_w;
            
            // CS goes low to start transaction (triggers snapshot)
            cs_n = 1'b0;
            #(5 * CLK_PERIOD);  // Setup time for first bit
            
            // Verify snapshot was captured
            $display("[%0t] MCU: Snapshot captured - quat1_w_snap=%d, quat1_w_input=%d", 
                     $time, quat1_w_snap, quat1_w);
            
            // Verify first bit is ready (should be MSB of 0xAA = 1)
            if (sdo == 1'b1) begin
                $display("[%0t] MCU: First bit ready (MSB=1) ✓", $time);
            end else begin
                $display("[%0t] MCU: ERROR - First bit not ready! sdo=%b", $time, sdo);
            end
            
            // Read 16 bytes (128 bits total)
            // SPI Mode 0: CPOL=0 (idle low), CPHA=0 (sample on rising, change on falling)
            for (i = 0; i < 16; i = i + 1) begin
                received_packet[i] = 8'h00;
                
                // Read 8 bits MSB first (SPI Mode 0: SCK starts low, first edge is rising)
                for (j = 7; j >= 0; j = j - 1) begin
                    // SPI Mode 0 timing:
                    // - Rising edge: MCU samples data
                    // - Falling edge: FPGA shifts to prepare next bit
                    
                    // Rising edge - MCU samples
                    sck = 1'b1;
                    #(10);  // Small delay for sampling
                    received_packet[i][j] = sdo;
                    #(SCK_PERIOD/2 - 10);
                    
                    // Debug output for first byte
                    if (i == 0 && j >= 4) begin
                        $display("[%0t] Bit %0d: sdo=%b, shift_out=0x%02X, bit_count=%0d", 
                                 $time, j, sdo, shift_out, bit_count);
                    end
                    
                    // Falling edge - FPGA shifts to prepare next bit (except after last bit)
                    if (j > 0 || i < 15) begin
                        sck = 1'b0;
                        #(SCK_PERIOD/2);
                    end
                end
                
                $display("[%0t] MCU: Byte[%0d] = 0x%02X", $time, i, received_packet[i]);
            end
            
            // Verify data stability: change input data during transaction
            // Snapshot should prevent this from affecting the transaction
            quat1_w = 16'hFFFF;  // Change input data
            #(CLK_PERIOD);
            
            // Verify snapshot data is still being used (not affected by input change)
            if (quat1_w_snap == data_before_transaction) begin
                $display("[%0t] MCU: Data stability verified - snapshot preserved", $time);
            end else begin
                $display("[%0t] MCU: WARNING - Snapshot may have changed!", $time);
            end
            
            // Restore original data
            quat1_w = data_before_transaction;
            
            // CS goes high to end transaction
            cs_n = 1'b1;
            #(5 * CLK_PERIOD);
            
            $display("[%0t] MCU: SPI transaction complete", $time);
        end
    endtask
    
    // Main test sequence
    initial begin
        $dumpfile("tb_spi_slave_mcu_debug.vcd");
        $dumpvars(0, tb_spi_slave_mcu_debug);
        
        $display("========================================");
        $display("MCU SPI Slave Debug Testbench");
        $display("========================================");
        $display("");
        
        // Initialize
        cs_n = 1'b1;  // CS high (idle)
        sck = 1'b0;   // SCK idle low (Mode 0)
        sdi = 1'b0;
        quat1_valid = 1'b1;
        gyro1_valid = 1'b1;
        
        // Set test data
        quat1_w = 16'h1234;
        quat1_x = 16'h5678;
        quat1_y = 16'h9ABC;
        quat1_z = 16'hDEF0;
        gyro1_x = 16'h1111;
        gyro1_y = 16'h2222;
        gyro1_z = 16'h3333;
        
        #(10 * CLK_PERIOD);
        
        // ========================================
        // TEST 1: Verify Packet Buffer Assembly
        // ========================================
        $display("=== Test 1: Packet Buffer Assembly ===");
        
        // Wait for combinational logic
        #(2 * CLK_PERIOD);
        
        // Check header
        check_test("Test 1.1: Header byte = 0xAA", 
                   dut.packet_buffer[0] == 8'hAA);
        
        // Check quaternion data
        check_test("Test 1.2: Quat W MSB/LSB", 
                   dut.packet_buffer[1] == 8'h12 && dut.packet_buffer[2] == 8'h34);
        check_test("Test 1.3: Quat X MSB/LSB", 
                   dut.packet_buffer[3] == 8'h56 && dut.packet_buffer[4] == 8'h78);
        
        // Check gyroscope data
        check_test("Test 1.4: Gyro X MSB/LSB", 
                   dut.packet_buffer[9] == 8'h11 && dut.packet_buffer[10] == 8'h11);
        
        // Check flags
        check_test("Test 1.5: Flags byte (both valid)", 
                   dut.packet_buffer[15] == 8'h03);
        
        $display("");
        
        // ========================================
        // TEST 2: CS Reset and First Byte Load
        // ========================================
        $display("=== Test 2: CS Reset and First Byte Load ===");
        
        // CS should be high initially
        check_test("Test 2.1: CS high initially", cs_n == 1'b1);
        
        // When CS goes high, shift_out should be loaded with first byte
        #(5 * CLK_PERIOD);
        check_test("Test 2.2: shift_out loaded when CS high", 
                   shift_out == 8'hAA);
        check_test("Test 2.3: byte_count reset when CS high", byte_count == 0);
        check_test("Test 2.4: bit_count reset when CS high", bit_count == 0);
        
        $display("");
        
        // ========================================
        // TEST 3: SPI Transaction - First Byte
        // ========================================
        $display("=== Test 3: SPI Transaction - First Byte (0xAA) ===");
        
        // CS goes low
        cs_n = 1'b0;
        #(5 * CLK_PERIOD);
        
        // First bit should be ready (MSB of 0xAA = 1)
        check_test("Test 3.1: First bit ready (MSB=1)", sdo == 1'b1);
        check_test("Test 3.2: shift_out still 0xAA", shift_out == 8'hAA);
        
        // Clock out first byte (SPI Mode 0: SCK starts low, first edge is rising)
        for (bit_idx = 7; bit_idx >= 0; bit_idx = bit_idx - 1) begin
            // Rising edge - MCU samples this bit
            sck = 1'b1;
            #(10);
            sampled_bit = sdo;
            #(SCK_PERIOD/2 - 10);
            
            // Verify bit value
            expected_bit = (8'hAA >> bit_idx) & 1'b1;
            check_test($sformatf("Test 3.3: Bit %0d = %b", bit_idx, expected_bit), 
                       sampled_bit == expected_bit);
            
            // Falling edge - FPGA shifts to prepare next bit (except after last bit)
            if (bit_idx > 0) begin
                sck = 1'b0;
                #(SCK_PERIOD/2);
            end
        end
        
        // SCK returns to idle low
        sck = 1'b0;
        #(SCK_PERIOD/2);
        
        // After 8 bits, byte_count should increment
        check_test("Test 3.4: byte_count incremented after first byte", 
                   byte_count == 1);
        check_test("Test 3.5: bit_count reset after first byte", bit_count == 0);
        
        $display("");
        
        // ========================================
        // TEST 4: Complete 16-Byte Transaction
        // ========================================
        $display("=== Test 4: Complete 16-Byte Transaction ===");
        
        // Reset CS and read complete packet
        cs_n = 1'b1;
        #(10 * CLK_PERIOD);
        
        mcu_read_packet_cs();
        
        // Verify header
        check_test("Test 4.1: Header byte = 0xAA", 
                   received_packet[0] == 8'hAA);
        
        // Verify quaternion data
        check_test("Test 4.2: Quat W = 0x1234", 
                   received_packet[1] == 8'h12 && received_packet[2] == 8'h34);
        check_test("Test 4.3: Quat X = 0x5678", 
                   received_packet[3] == 8'h56 && received_packet[4] == 8'h78);
        
        // Verify gyroscope data
        check_test("Test 4.4: Gyro X = 0x1111", 
                   received_packet[9] == 8'h11 && received_packet[10] == 8'h11);
        
        // Verify flags
        check_test("Test 4.5: Flags = 0x03", 
                   received_packet[15] == 8'h03);
        
        $display("");
        
        // ========================================
        // TEST 5: Data Stability During Transaction
        // ========================================
        $display("=== Test 5: Data Stability During Transaction ===");
        
        // Reset
        cs_n = 1'b1;
        #(10 * CLK_PERIOD);
        
        // Set initial data
        quat1_w = 16'hABCD;
        quat1_x = 16'h1234;
        #(10 * CLK_PERIOD);
        
        // Start transaction
        cs_n = 1'b0;
        #(5 * CLK_PERIOD);
        
        // Verify snapshot was captured
        check_test("Test 5.1: Snapshot captured quat1_w", quat1_w_snap == 16'hABCD);
        check_test("Test 5.2: Snapshot captured quat1_x", quat1_x_snap == 16'h1234);
        
        // Change input data during transaction (should not affect snapshot)
        quat1_w = 16'hFFFF;
        quat1_x = 16'h0000;
        #(CLK_PERIOD);
        
        // Verify snapshot is unchanged
        check_test("Test 5.3: Snapshot preserved during transaction (quat1_w)", 
                   quat1_w_snap == 16'hABCD);
        check_test("Test 5.4: Snapshot preserved during transaction (quat1_x)", 
                   quat1_x_snap == 16'h1234);
        
        // Read a few bytes to verify data is from snapshot
        for (i = 0; i < 2; i = i + 1) begin
            for (j = 7; j >= 0; j = j - 1) begin
                // Rising edge - MCU samples
                sck = 1'b1;
                #(SCK_PERIOD/2);
                // Falling edge - FPGA shifts
                sck = 1'b0;
                #(SCK_PERIOD/2);
            end
        end
        
        // Verify snapshot still unchanged
        check_test("Test 5.5: Snapshot still preserved after partial read", 
                   quat1_w_snap == 16'hABCD);
        
        cs_n = 1'b1;
        #(10 * CLK_PERIOD);
        
        $display("");
        
        // ========================================
        // TEST 6: Clock Domain Crossing Verification
        // ========================================
        $display("=== Test 6: Clock Domain Crossing ===");
        
        // Set data in clk domain
        quat1_w = 16'h5678;
        quat1_valid = 1'b1;
        #(10 * CLK_PERIOD);  // Allow data to propagate in clk domain
        
        // CS falling edge should capture synchronized data
        cs_n = 1'b0;
        #(5 * CLK_PERIOD);
        
        // Verify snapshot captured the data (may have slight delay due to CDC)
        // Allow some time for synchronization
        #(2 * CLK_PERIOD);
        check_test("Test 6.1: Snapshot captured data after CDC", 
                   quat1_w_snap == 16'h5678 || quat1_w_snap == 16'h0000);  // May be 0 if not synced yet
        
        cs_n = 1'b1;
        #(10 * CLK_PERIOD);
        
        $display("");
        
        // ========================================
        // Summary
        // ========================================
        $display("========================================");
        $display("Test Summary");
        $display("========================================");
        $display("Total Tests: %0d", test_count);
        $display("Passed: %0d", pass_count);
        $display("Failed: %0d", fail_count);
        $display("========================================");
        
        if (fail_count == 0) begin
            $display("ALL TESTS PASSED");
        end else begin
            $display("SOME TESTS FAILED");
        end
        $display("========================================");
        
        #(100 * CLK_PERIOD);
        $finish;
    end
    
endmodule


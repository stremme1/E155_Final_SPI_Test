// Sadhvi Narayanan, sanarayanan@g.hmc.edu, 10/26/2025
// aes spi module to handle spi transactions with the FPGA

/////////////////////////////////////////////
// aes_spi
//   SPI interface.  Shifts in key and plaintext
//   Captures ciphertext when done, then shifts it out
//   Tricky cases to properly change sdo on negedge clk
/////////////////////////////////////////////
module aes_spi(input  logic sck,
             input  logic sdi,
             output logic sdo,
             input  logic done,
             output logic [127:0] key, plaintext,
             input  logic [127:0] cyphertext);


  logic         sdodelayed, wasdone;
  logic [127:0] cyphertextcaptured;
           
  // assert load
  // apply 256 sclks to shift in key and plaintext, starting with plaintext[127]
  // then deassert load, wait until done
  // then apply 128 sclks to shift out cyphertext, starting with cyphertext[127]
  // SPI mode is equivalent to cpol = 0, cpha = 0 since data is sampled on first edge and the first
  // edge is a rising edge (clock going from low in the idle state to high).
  always_ff @(posedge sck)
      if (!wasdone)  {cyphertextcaptured, plaintext, key} = {cyphertext, plaintext[126:0], key, sdi};
      else           {cyphertextcaptured, plaintext, key} = {cyphertextcaptured[126:0], plaintext, key, sdi};
   // sdo should change on the negative edge of sck
  always_ff @(negedge sck) begin
      wasdone = done;
      sdodelayed = cyphertextcaptured[126];
  end
   // when done is first asserted, shift out msb before clock edge
  assign sdo = (done & !wasdone) ? cyphertext[127] : sdodelayed;
endmodule
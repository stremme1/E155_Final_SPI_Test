`timescale 1ns / 1ps

// Testbench for Arduino SPI Slave Module
// Tests SPI slave operation for receiving 16-byte packets from Arduino
// Verifies packet reception, header validation, and data mapping to MCU interface
// SPI Mode 0 (CPOL=0, CPHA=0) at 100kHz (10us period)

module tb_arduino_spi_slave;

    // Clock
    logic clk;
    
    // Arduino SPI interface (Arduino is master, FPGA is slave)
    logic cs_n;      // Chip select from Arduino (active low)
    logic sck;       // SPI clock from Arduino
    logic sdi;       // SPI data in (MOSI from Arduino)
    
    // DUT outputs
    logic initialized;
    logic error;
    logic quat1_valid;
    logic signed [15:0] quat1_w, quat1_x, quat1_y, quat1_z;
    logic gyro1_valid;
    logic signed [15:0] gyro1_x, gyro1_y, gyro1_z;
    
    // Clock generation (3MHz FPGA clock)
    parameter CLK_PERIOD = 333;  // 3MHz = 333ns period
    always begin
        clk = 0;
        #(CLK_PERIOD/2);
        clk = 1;
        #(CLK_PERIOD/2);
    end
    
    // Arduino SPI clock - 100kHz (10us period = 10000ns)
    // SCK starts idle low (SPI Mode 0: CPOL=0)
    parameter SCK_PERIOD = 10000;  // 100kHz = 10us period
    initial begin
        sck = 0;  // Idle low for SPI Mode 0
    end
    
    // DUT
    arduino_spi_slave dut (
        .clk(clk),
        .cs_n(cs_n),
        .sck(sck),
        .sdi(sdi),
        .initialized(initialized),
        .error(error),
        .quat1_valid(quat1_valid),
        .quat1_w(quat1_w),
        .quat1_x(quat1_x),
        .quat1_y(quat1_y),
        .quat1_z(quat1_z),
        .gyro1_valid(gyro1_valid),
        .gyro1_x(gyro1_x),
        .gyro1_y(gyro1_y),
        .gyro1_z(gyro1_z)
    );
    
    // Access internal signals for debugging
    wire [7:0] packet_buffer_0 = dut.packet_buffer[0];
    wire [7:0] packet_buffer_1 = dut.packet_buffer[1];
    wire [7:0] packet_buffer_2 = dut.packet_buffer[2];
    wire [3:0] byte_count = dut.byte_count;
    wire [2:0] bit_count = dut.bit_count;
    wire [7:0] rx_shift = dut.rx_shift;
    wire [7:0] header = dut.header;
    wire signed [15:0] roll = dut.roll;
    wire signed [15:0] pitch = dut.pitch;
    wire signed [15:0] yaw = dut.yaw;
    
    // Test tracking
    integer test_count = 0;
    integer pass_count = 0;
    integer fail_count = 0;
    
    // Helper task to check and report
    task check_test(input string test_name, input logic condition);
        test_count = test_count + 1;
        if (condition) begin
            $display("[PASS] %s", test_name);
            pass_count = pass_count + 1;
        end else begin
            $display("[FAIL] %s", test_name);
            fail_count = fail_count + 1;
        end
    endtask
    
    // Helper task to wait for clock domain crossing
    task wait_cdc;
        #(CLK_PERIOD * 20);  // Wait 20 clock cycles for CDC and packet processing
    endtask
    
    // Task to send a byte via SPI (MSB first, Mode 0)
    // Assumes CS is already low
    // For MSB-first: send bit 7 first, then bit 6, ..., then bit 0
    task send_spi_byte(input [7:0] data);
        integer i;
        $display("    [SPI] Sending byte: 0x%02X (binary: %b)", data, data);
        for (i = 7; i >= 0; i = i - 1) begin
            // Set data before rising edge (setup time)
            sdi = data[i];
            #(SCK_PERIOD/4);  // Setup time
            sck = 1;  // Rising edge - FPGA samples sdi here
            #(SCK_PERIOD/4);  // Hold time
            // $display("      Bit %0d: sdi=%b (from data[%0d]=%b)", 7-i, sdi, i, data[i]);
            #(SCK_PERIOD/2);
            sck = 0;  // Falling edge
        end
        $display("    [SPI] Byte sent: 0x%02X", data);
    endtask
    
    // Task to send a complete 16-byte packet (inline version to avoid unpacked array issues)
    task send_packet_inline;
        input [7:0] b0, b1, b2, b3, b4, b5, b6, b7, b8, b9, b10, b11, b12, b13, b14, b15;
        // CS falling edge - ensure CS is high first, then go low
        cs_n = 1;
        #(SCK_PERIOD * 3);  // Wait longer to ensure CS is stable high
        cs_n = 0;
        #(SCK_PERIOD * 2);  // Wait for CS to stabilize low before first SCK edge
        
        // Send all 16 bytes
        send_spi_byte(b0);
        send_spi_byte(b1);
        send_spi_byte(b2);
        send_spi_byte(b3);
        send_spi_byte(b4);
        send_spi_byte(b5);
        send_spi_byte(b6);
        send_spi_byte(b7);
        send_spi_byte(b8);
        send_spi_byte(b9);
        send_spi_byte(b10);
        send_spi_byte(b11);
        send_spi_byte(b12);
        send_spi_byte(b13);
        send_spi_byte(b14);
        send_spi_byte(b15);
        
        // CS rising edge (transaction complete)
        #(SCK_PERIOD);
        cs_n = 1;
        #(SCK_PERIOD * 3);  // Wait longer for CS to stabilize high
    endtask
    
    // Main test sequence
    initial begin
        $dumpfile("tb_arduino_spi_slave.vcd");
        $dumpvars(0, tb_arduino_spi_slave);
        
        $display("========================================");
        $display("Arduino SPI Slave Testbench");
        $display("========================================");
        $display("");
        
        // Initialize
        cs_n = 1;
        sck = 0;
        sdi = 0;
        
        #(10 * CLK_PERIOD);
        
        // ========================================
        // TEST 0: Bit Shifting Verification
        // ========================================
        $display("=== Test 0: Bit Shifting Verification ===");
        
        // Test 0.1: Send 0xAA to verify MSB-first bit order
        begin
            $display("Test 0.1: Sending 0xAA to verify bit shifting");
            cs_n = 1;
            #(SCK_PERIOD * 3);
            cs_n = 0;
            #(SCK_PERIOD * 2);
            
            send_spi_byte(8'hAA);  // 0xAA = 0b10101010
            
            // CS rising edge
            #(SCK_PERIOD);
            cs_n = 1;
            #(SCK_PERIOD * 3);
            
            // Wait for CDC
            wait(cs_n == 1'b1);
            repeat(20) @(posedge clk);
            
            // Check if byte was received correctly
            $display("    packet_buffer[0] = 0x%02X (expected 0xAA)", packet_buffer_0);
            check_test("Test 0.1: Byte 0xAA received correctly", packet_buffer_0 == 8'hAA);
            $display("    Expected: First bit=1 (MSB), Last bit=0 (LSB)");
            $display("    Pattern: 1-0-1-0-1-0-1-0");
        end
        
        // Test 0.2: Send 0x55 to verify opposite pattern
        begin
            $display("Test 0.2: Sending 0x55 to verify bit shifting");
            cs_n = 1;
            #(SCK_PERIOD * 3);
            cs_n = 0;
            #(SCK_PERIOD * 2);
            
            send_spi_byte(8'h55);  // 0x55 = 0b01010101
            
            // CS rising edge
            #(SCK_PERIOD);
            cs_n = 1;
            #(SCK_PERIOD * 3);
            
            // Wait for CDC
            wait(cs_n == 1'b1);
            repeat(20) @(posedge clk);
            
            $display("    packet_buffer[0] = 0x%02X (expected 0x55)", packet_buffer_0);
            check_test("Test 0.2: Byte 0x55 received correctly", packet_buffer_0 == 8'h55);
            $display("    Expected: First bit=0 (MSB), Last bit=1 (LSB)");
            $display("    Pattern: 0-1-0-1-0-1-0-1");
        end
        
        $display("");
        
        // ========================================
        // TEST 1: Valid Packet Reception
        // ========================================
        $display("=== Test 1: Valid Packet Reception ===");
        
        // Test 1.1: Valid packet with header 0xAA
        begin
            $display("Test 1.1: Sending valid packet with header 0xAA");
            // Header = 0xAA
            // Roll = 1000 (0.01° resolution = 10.00°)
            // Pitch = -500 (-5.00°)
            // Yaw = 2000 (20.00°)
            // Gyro X = 100, Y = -200, Z = 50
            // Flags: both valid (0x03)
            send_packet_inline(
                8'hAA,  // Header
                8'h03, 8'hE8,  // Roll = 1000
                8'hFE, 8'h0C,  // Pitch = -500
                8'h07, 8'hD0,  // Yaw = 2000
                8'h00, 8'h64,  // Gyro X = 100
                8'hFF, 8'h38,  // Gyro Y = -200
                8'h00, 8'h32,  // Gyro Z = 50
                8'h03,  // Flags: both valid
                8'h00, 8'h00   // Reserved
            );
            // Wait for CS rising edge to be detected and packet to be processed
            // Wait for CS to go high, then wait for synchronization and processing
            wait(cs_n == 1'b1);  // Wait for CS to go high
            repeat(25) @(posedge clk);  // Wait for CDC synchronization (increased for stability)
            
            // Debug output - check internal signals
            $display("    Internal signals after packet reception:");
            $display("      packet_buffer[0] = 0x%02X (header, expected 0xAA)", packet_buffer_0);
            $display("      packet_buffer[1] = 0x%02X (Roll MSB, expected 0x03)", packet_buffer_1);
            $display("      packet_buffer[2] = 0x%02X (Roll LSB, expected 0xE8)", packet_buffer_2);
            $display("      header = 0x%02X, roll = 0x%04X (%0d)", header, roll, roll);
            $display("      pitch = 0x%04X (%0d), yaw = 0x%04X (%0d)", pitch, pitch, yaw, yaw);
            
            // Debug output - check outputs
            $display("    Output signals after packet reception:");
            $display("      initialized = %b, error = %b", initialized, error);
            $display("      quat1_w = 0x%04X (%0d), quat1_x = 0x%04X (%0d)", quat1_w, quat1_w, quat1_x, quat1_x);
            $display("      quat1_y = 0x%04X (%0d), quat1_z = 0x%04X (%0d)", quat1_y, quat1_y, quat1_z, quat1_z);
            $display("      gyro1_x = 0x%04X (%0d), gyro1_y = 0x%04X (%0d), gyro1_z = 0x%04X (%0d)", 
                     gyro1_x, gyro1_x, gyro1_y, gyro1_y, gyro1_z, gyro1_z);
            $display("      quat1_valid = %b, gyro1_valid = %b", quat1_valid, gyro1_valid);
            
            // Check outputs
            check_test("Test 1.1a: Header valid → initialized = 1", initialized == 1'b1);
            check_test("Test 1.1b: Header valid → error = 0", error == 1'b0);
            check_test("Test 1.1c: Quat W = 16384 (Q14 format)", quat1_w == 16'd16384);
            check_test("Test 1.1d: Quat X = Roll (1000)", quat1_x == 16'd1000);
            check_test("Test 1.1e: Quat Y = Pitch (-500)", quat1_y == -16'd500);
            check_test("Test 1.1f: Quat Z = Yaw (2000)", quat1_z == 16'd2000);
            check_test("Test 1.1g: Gyro X = 100", gyro1_x == 16'd100);
            check_test("Test 1.1h: Gyro Y = -200", gyro1_y == -16'd200);
            check_test("Test 1.1i: Gyro Z = 50", gyro1_z == 16'd50);
            check_test("Test 1.1j: Quat valid = 1 (from flags[0])", quat1_valid == 1'b1);
            check_test("Test 1.1k: Gyro valid = 1 (from flags[1])", gyro1_valid == 1'b1);
        end
        
        $display("");
        
        // ========================================
        // TEST 2: Invalid Header Detection
        // ========================================
        $display("=== Test 2: Invalid Header Detection ===");
        
        // Test 2.1: Invalid header (0x55 instead of 0xAA)
        begin
            send_packet_inline(
                8'h55,  // Invalid header
                8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,  // Roll, Pitch, Yaw
                8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,  // Gyro X, Y, Z
                8'h00,  // Flags
                8'h00, 8'h00   // Reserved
            );
            wait_cdc();
            
            check_test("Test 2.1a: Invalid header → initialized = 0", initialized == 1'b0);
            check_test("Test 2.1b: Invalid header → error = 1", error == 1'b1);
        end
        
        // Test 2.2: Valid header restores status
        begin
            send_packet_inline(
                8'hAA,  // Valid header
                8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,  // Roll, Pitch, Yaw
                8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,  // Gyro X, Y, Z
                8'h03,  // Flags: both valid
                8'h00, 8'h00   // Reserved
            );
            wait_cdc();
            
            check_test("Test 2.2a: Valid header restores initialized = 1", initialized == 1'b1);
            check_test("Test 2.2b: Valid header clears error = 0", error == 1'b0);
        end
        
        $display("");
        
        // ========================================
        // TEST 3: Flag Mapping
        // ========================================
        $display("=== Test 3: Flag Mapping ===");
        
        // Test 3.1: Only Euler valid (flag = 0x01)
        begin
            send_packet_inline(
                8'hAA,  // Header
                8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,  // Roll, Pitch, Yaw
                8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,  // Gyro X, Y, Z
                8'h01,  // Flags: only Euler valid
                8'h00, 8'h00   // Reserved
            );
            wait_cdc();
            
            check_test("Test 3.1a: Flag 0x01 → quat_valid = 1", quat1_valid == 1'b1);
            check_test("Test 3.1b: Flag 0x01 → gyro_valid = 0", gyro1_valid == 1'b0);
        end
        
        // Test 3.2: Only Gyro valid (flag = 0x02)
        begin
            send_packet_inline(
                8'hAA,  // Header
                8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,  // Roll, Pitch, Yaw
                8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,  // Gyro X, Y, Z
                8'h02,  // Flags: only Gyro valid
                8'h00, 8'h00   // Reserved
            );
            wait_cdc();
            
            check_test("Test 3.2a: Flag 0x02 → quat_valid = 0", quat1_valid == 1'b0);
            check_test("Test 3.2b: Flag 0x02 → gyro_valid = 1", gyro1_valid == 1'b1);
        end
        
        // Test 3.3: Both valid (flag = 0x03)
        begin
            send_packet_inline(
                8'hAA,  // Header
                8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,  // Roll, Pitch, Yaw
                8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,  // Gyro X, Y, Z
                8'h03,  // Flags: both valid
                8'h00, 8'h00   // Reserved
            );
            wait_cdc();
            
            check_test("Test 3.3a: Flag 0x03 → quat_valid = 1", quat1_valid == 1'b1);
            check_test("Test 3.3b: Flag 0x03 → gyro_valid = 1", gyro1_valid == 1'b1);
        end
        
        // Test 3.4: Neither valid (flag = 0x00)
        begin
            send_packet_inline(
                8'hAA,  // Header
                8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,  // Roll, Pitch, Yaw
                8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,  // Gyro X, Y, Z
                8'h00,  // Flags: neither valid
                8'h00, 8'h00   // Reserved
            );
            wait_cdc();
            
            check_test("Test 3.4a: Flag 0x00 → quat_valid = 0", quat1_valid == 1'b0);
            check_test("Test 3.4b: Flag 0x00 → gyro_valid = 0", gyro1_valid == 1'b0);
        end
        
        $display("");
        
        // ========================================
        // TEST 4: Edge Cases
        // ========================================
        $display("=== Test 4: Edge Cases ===");
        
        // Test 4.1: Maximum positive values
        begin
            send_packet_inline(
                8'hAA,  // Header
                8'h7F, 8'hFF,  // Roll = 32767
                8'h7F, 8'hFF,  // Pitch = 32767
                8'h7F, 8'hFF,  // Yaw = 32767
                8'h7F, 8'hFF,  // Gyro X = 32767
                8'h7F, 8'hFF,  // Gyro Y = 32767
                8'h7F, 8'hFF,  // Gyro Z = 32767
                8'h03,  // Flags: both valid
                8'h00, 8'h00   // Reserved
            );
            wait_cdc();
            
            check_test("Test 4.1a: Max positive Roll (32767)", quat1_x == 16'd32767);
            check_test("Test 4.1b: Max positive Pitch (32767)", quat1_y == 16'd32767);
            check_test("Test 4.1c: Max positive Yaw (32767)", quat1_z == 16'd32767);
            check_test("Test 4.1d: Max positive Gyro X (32767)", gyro1_x == 16'd32767);
        end
        
        // Test 4.2: Maximum negative values
        begin
            send_packet_inline(
                8'hAA,  // Header
                8'h80, 8'h00,  // Roll = -32768
                8'h80, 8'h00,  // Pitch = -32768
                8'h80, 8'h00,  // Yaw = -32768
                8'h80, 8'h00,  // Gyro X = -32768
                8'h80, 8'h00,  // Gyro Y = -32768
                8'h80, 8'h00,  // Gyro Z = -32768
                8'h03,  // Flags: both valid
                8'h00, 8'h00   // Reserved
            );
            wait_cdc();
            
            check_test("Test 4.2a: Max negative Roll (-32768)", quat1_x == -16'd32768);
            check_test("Test 4.2b: Max negative Pitch (-32768)", quat1_y == -16'd32768);
            check_test("Test 4.2c: Max negative Yaw (-32768)", quat1_z == -16'd32768);
            check_test("Test 4.2d: Max negative Gyro X (-32768)", gyro1_x == -16'd32768);
        end
        
        // Test 4.3: Zero values
        begin
            send_packet_inline(
                8'hAA,  // Header
                8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,  // Roll, Pitch, Yaw = 0
                8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,  // Gyro X, Y, Z = 0
                8'h03,  // Flags: both valid
                8'h00, 8'h00   // Reserved
            );
            wait_cdc();
            
            check_test("Test 4.3a: Zero Roll", quat1_x == 16'd0);
            check_test("Test 4.3b: Zero Pitch", quat1_y == 16'd0);
            check_test("Test 4.3c: Zero Yaw", quat1_z == 16'd0);
            check_test("Test 4.3d: Zero Gyro X", gyro1_x == 16'd0);
        end
        
        $display("");
        
        // ========================================
        // TEST 5: Multiple Packets
        // ========================================
        $display("=== Test 5: Multiple Packets ===");
        
        // Test 5.1: Send multiple packets and verify data updates
        begin
            // First packet: Roll = 100
            send_packet_inline(
                8'hAA,  // Header
                8'h00, 8'h64,  // Roll = 100
                8'h00, 8'h00,  // Pitch = 0
                8'h00, 8'h00,  // Yaw = 0
                8'h00, 8'h00,  // Gyro X = 0
                8'h00, 8'h00,  // Gyro Y = 0
                8'h00, 8'h00,  // Gyro Z = 0
                8'h03,  // Flags: both valid
                8'h00, 8'h00   // Reserved
            );
            wait_cdc();
            check_test("Test 5.1a: First packet Roll = 100", quat1_x == 16'd100);
            
            // Second packet: Roll = 500
            send_packet_inline(
                8'hAA,  // Header
                8'h01, 8'hF4,  // Roll = 500
                8'h00, 8'h00,  // Pitch = 0
                8'h00, 8'h00,  // Yaw = 0
                8'h00, 8'h00,  // Gyro X = 0
                8'h00, 8'h00,  // Gyro Y = 0
                8'h00, 8'h00,  // Gyro Z = 0
                8'h03,  // Flags: both valid
                8'h00, 8'h00   // Reserved
            );
            wait_cdc();
            check_test("Test 5.1b: Second packet Roll = 500", quat1_x == 16'd500);
        end
        
        $display("");
        
        // ========================================
        // Summary
        // ========================================
        $display("========================================");
        $display("Test Summary");
        $display("========================================");
        $display("Total Tests: %0d", test_count);
        $display("Passed: %0d", pass_count);
        $display("Failed: %0d", fail_count);
        $display("========================================");
        
        if (fail_count == 0) begin
            $display("ALL TESTS PASSED");
        end else begin
            $display("SOME TESTS FAILED");
        end
        $display("========================================");
        
        #(10 * CLK_PERIOD);
        $finish;
    end
    
endmodule


`timescale 1ns / 1ps

// MCU SPI Slave Module
// FPGA is SPI slave to MCU (MCU is master) - READ-ONLY MODE
// Sends RAW sensor data packets to MCU
// Based on e155-lab7-main 2/fpga/src/aes_spi.sv pattern
// SPI Mode 0 (CPOL=0, CPHA=0): MCU samples on rising edge, FPGA changes on falling edge
// 
// Read-Only Protocol:
// - FPGA ignores MOSI (sdi) completely - only shifts out data on MISO (sdo)
// - MCU generates SCK by sending dummy bytes (0x00) via spiSendReceive(0)
// - FPGA shifts out 1 bit per SCK edge from its shift register
// - MCU reads data from MISO during the transaction

module spi_slave_mcu(
    input  logic        clk,           // FPGA system clock
    input  logic        sck,           // SPI clock from MCU (generated by MCU)
    input  logic        sdi,           // SPI data in (MOSI from MCU - IGNORED in read-only mode)
    output logic        sdo,           // SPI data out (MISO to MCU - shifts out data)
    input  logic        load,          // Load signal from MCU (acknowledge)
    output logic        done,          // Done signal to MCU (data ready)
    
    // Sensor data inputs (RAW data from BNO085 controller)
    // Sensor 1 (Right Hand) - Single sensor only
    input  logic        quat1_valid,
    input  logic signed [15:0] quat1_w, quat1_x, quat1_y, quat1_z,
    input  logic        gyro1_valid,
    input  logic signed [15:0] gyro1_x, gyro1_y, gyro1_z
);

    // Packet format: 16 bytes total (single sensor only)
    // Byte 0:    Header (0xAA)
    // Byte 1-8:  Sensor 1 Quaternion (w, x, y, z - MSB,LSB each)
    // Byte 9-14: Sensor 1 Gyroscope (x, y, z - MSB,LSB each)
    // Byte 15:   Sensor 1 Flags (bit 0=quat_valid, bit 1=gyro_valid)
    
    localparam PACKET_SIZE = 16;
    localparam HEADER_BYTE = 8'hAA;
    
    // Packet buffer - assembled from sensor data
    logic [7:0] packet_buffer [0:PACKET_SIZE-1];
    logic [7:0] tx_shift_reg;
    logic       sdodelayed, wasdone;
    logic       data_ready;
    logic       load_prev;
    logic [4:0] bit_cnt;  // 5 bits for 16 bytes * 8 bits = 128 bits
    
    // Assemble packet from sensor data (using assign statements for iverilog compatibility)
    // Header
    assign packet_buffer[0] = HEADER_BYTE;
    
    // Sensor 1 Quaternion (MSB,LSB format)
    assign packet_buffer[1] = quat1_w[15:8];  // W MSB
    assign packet_buffer[2] = quat1_w[7:0];   // W LSB
    assign packet_buffer[3] = quat1_x[15:8];  // X MSB
    assign packet_buffer[4] = quat1_x[7:0];   // X LSB
    assign packet_buffer[5] = quat1_y[15:8];  // Y MSB
    assign packet_buffer[6] = quat1_y[7:0];   // Y LSB
    assign packet_buffer[7] = quat1_z[15:8];  // Z MSB
    assign packet_buffer[8] = quat1_z[7:0];   // Z LSB
    
    // Sensor 1 Gyroscope (MSB,LSB format)
    assign packet_buffer[9]  = gyro1_x[15:8];  // X MSB
    assign packet_buffer[10] = gyro1_x[7:0];   // X LSB
    assign packet_buffer[11] = gyro1_y[15:8];  // Y MSB
    assign packet_buffer[12] = gyro1_y[7:0];   // Y LSB
    assign packet_buffer[13] = gyro1_z[15:8];  // Z MSB
    assign packet_buffer[14] = gyro1_z[7:0];   // Z LSB
    
    // Sensor 1 Flags
    assign packet_buffer[15] = {6'h0, gyro1_valid, quat1_valid};
    
    // Data ready when either sensor has valid data
    // Simplified logic: detect 0->1 transition on has_valid, clear on LOAD acknowledgment
    logic data_ready_reg = 1'b0;
    logic has_valid;
    logic has_valid_prev = 1'b0;
    logic load_prev = 1'b0;
    
    // TEST MODE: Force DONE to assert after a delay (for testing SPI communication)
    // Set to 1 to enable test mode, 0 for normal operation
    localparam TEST_MODE = 1'b0;  // Change to 1'b1 to force DONE assertion
    logic [23:0] init_delay_counter = 24'd0;
    logic test_done = 1'b0;
    
    assign has_valid = (quat1_valid || gyro1_valid);
    
    always_ff @(posedge clk) begin
        load_prev <= load;
        
        // TEST MODE: Force DONE after initialization delay
        if (TEST_MODE) begin
            if (init_delay_counter < 24'd3_000_000) begin  // ~1 second @ 3MHz
                init_delay_counter <= init_delay_counter + 1;
                test_done <= 1'b0;
            end else begin
                test_done <= 1'b1;  // Force DONE high for testing
            end
        end else begin
            test_done <= 1'b0;
        end
        
        // Check for LOAD edge (acknowledgment) - highest priority
        if (load && !load_prev) begin
            // MCU acknowledged - clear data ready
            data_ready_reg <= 1'b0;
            has_valid_prev <= 1'b0;
        end else if (!TEST_MODE) begin
            // If valid data is present and we haven't seen it before, set data ready
            // This captures the one-cycle pulse from the BNO085 controller
            if (has_valid && !has_valid_prev) begin
                // New valid data detected - set data ready
                data_ready_reg <= 1'b1;
                has_valid_prev <= 1'b1;
            end else if (!has_valid) begin
                // No valid data - update tracking but keep data_ready_reg set
                // (it will be cleared by LOAD acknowledgment)
                has_valid_prev <= 1'b0;
            end
            // If has_valid && has_valid_prev, keep data_ready_reg set (already asserted)
        end
    end
    
    // Done signal: Assert when data is ready (or in test mode)
    assign done = TEST_MODE ? test_done : data_ready_reg;
    
    // Create a 128-bit shift register from packet buffer (16 bytes * 8 bits)
    // Read-only mode: FPGA ignores MOSI (sdi), only shifts out data on MISO (sdo)
    logic [127:0] packet_shift_reg;
    
    // SPI Mode 0 (CPOL=0, CPHA=0): MCU samples on rising edge, FPGA changes on falling edge
    // Shift register behavior:
    // - On first posedge when data ready: load packet_buffer into shift register (MSB first)
    // - On subsequent posedges: shift left (MSB first) - FPGA ignores SDI (MOSI)
    // - On negedge: update output for next bit
    always_ff @(posedge sck) begin
        if (!wasdone) begin
            // First posedge: load packet buffer into shift register (MSB first)
            // Pack all bytes: packet_buffer[0] is MSB of first byte, goes to bit 127
            // Read-only mode: ignore SDI (MOSI), only shift out data
            packet_shift_reg = {
                packet_buffer[0], packet_buffer[1], packet_buffer[2], packet_buffer[3],
                packet_buffer[4], packet_buffer[5], packet_buffer[6], packet_buffer[7],
                packet_buffer[8], packet_buffer[9], packet_buffer[10], packet_buffer[11],
                packet_buffer[12], packet_buffer[13], packet_buffer[14], packet_buffer[15]
            };
        end else begin
            // Subsequent posedges: shift left (MSB first)
            // Read-only mode: ignore SDI, shift in 0 (or just shift left)
            packet_shift_reg = {packet_shift_reg[126:0], 1'b0};
        end
    end
    
    // Track previous done state (for edge detection)
    // Update output on negedge (when FPGA should change MISO for next bit)
    // SPI Mode 0: FPGA changes MISO on falling edge, MCU samples on rising edge
    always_ff @(negedge sck) begin
        wasdone = done;  // Blocking assignment for immediate update
        // After shift on posedge, next bit to output is at bit 126 (was at 127 before shift)
        sdodelayed = packet_shift_reg[126];  // Next bit to output (MSB of remaining data)
    end
    
    // SDO (MISO) output: Read-only mode
    // SPI Mode 0 timing:
    // - Before first posedge: output MSB directly (done & !wasdone) = packet_buffer[0][7]
    // - After first negedge: wasdone becomes true, use sdodelayed (set on negedge)
    // packet_buffer[0][7] is MSB of first byte (bit 7 of byte 0), which is MSB of entire packet
    // sdodelayed is updated on negedge to packet_shift_reg[126] (next bit after shift)
    assign sdo = (done & !wasdone) ? packet_buffer[0][7] : sdodelayed;
    
endmodule



`timescale 1ns / 1ps

// MCU SPI Slave Module
// FPGA is SPI slave to MCU (MCU is master)
// Sends RAW sensor data packets to MCU
// Based on e155-lab7-main 2/fpga/src/aes_spi.sv pattern
// SPI Mode 0 (CPOL=0, CPHA=0): data sampled on rising edge, changed on falling edge

module mcu_spi_slave(
    input  logic        clk,           // FPGA system clock
    input  logic        sck,           // SPI clock from MCU
    input  logic        sdi,           // SPI data in (MOSI from MCU, not used for commands)
    output logic        sdo,           // SPI data out (MISO to MCU)
    input  logic        load,          // Load signal from MCU (acknowledge)
    output logic        done,          // Done signal to MCU (data ready)
    
    // Sensor data inputs (RAW data from BNO085 controllers)
    // Sensor 1 (Right Hand)
    input  logic        quat1_valid,
    input  logic signed [15:0] quat1_w, quat1_x, quat1_y, quat1_z,
    input  logic        gyro1_valid,
    input  logic signed [15:0] gyro1_x, gyro1_y, gyro1_z,
    
    // Sensor 2 (Left Hand)
    input  logic        quat2_valid,
    input  logic signed [15:0] quat2_w, quat2_x, quat2_y, quat2_z,
    input  logic        gyro2_valid,
    input  logic signed [15:0] gyro2_x, gyro2_y, gyro2_z
);

    // Packet format: 32 bytes total
    // Byte 0:    Header (0xAA)
    // Byte 1-8:  Sensor 1 Quaternion (w, x, y, z - MSB,LSB each)
    // Byte 9-14: Sensor 1 Gyroscope (x, y, z - MSB,LSB each)
    // Byte 15:   Sensor 1 Flags (bit 0=quat_valid, bit 1=gyro_valid)
    // Byte 16-23: Sensor 2 Quaternion (w, x, y, z - MSB,LSB each)
    // Byte 24-29: Sensor 2 Gyroscope (x, y, z - MSB,LSB each)
    // Byte 30:   Sensor 2 Flags (bit 0=quat_valid, bit 1=gyro_valid)
    // Byte 31:   Reserved (0x00)
    
    localparam PACKET_SIZE = 32;
    localparam HEADER_BYTE = 8'hAA;
    
    // Packet buffer - assembled from sensor data
    logic [7:0] packet_buffer [0:PACKET_SIZE-1];
    logic [7:0] tx_shift_reg;
    logic       sdodelayed, wasdone;
    logic       data_ready;
    logic       load_prev;
    logic [5:0] bit_cnt;  // 6 bits for 32 bytes * 8 bits = 256 bits
    
    // Assemble packet from sensor data (update continuously as data changes)
    always_comb begin
        // Header
        packet_buffer[0] = HEADER_BYTE;
        
        // Sensor 1 Quaternion (MSB,LSB format)
        packet_buffer[1] = quat1_w[15:8];  // W MSB
        packet_buffer[2] = quat1_w[7:0];   // W LSB
        packet_buffer[3] = quat1_x[15:8];  // X MSB
        packet_buffer[4] = quat1_x[7:0];   // X LSB
        packet_buffer[5] = quat1_y[15:8];  // Y MSB
        packet_buffer[6] = quat1_y[7:0];   // Y LSB
        packet_buffer[7] = quat1_z[15:8];  // Z MSB
        packet_buffer[8] = quat1_z[7:0];   // Z LSB
        
        // Sensor 1 Gyroscope (MSB,LSB format)
        packet_buffer[9]  = gyro1_x[15:8];  // X MSB
        packet_buffer[10] = gyro1_x[7:0];   // X LSB
        packet_buffer[11] = gyro1_y[15:8];  // Y MSB
        packet_buffer[12] = gyro1_y[7:0];   // Y LSB
        packet_buffer[13] = gyro1_z[15:8];  // Z MSB
        packet_buffer[14] = gyro1_z[7:0];   // Z LSB
        
        // Sensor 1 Flags
        packet_buffer[15] = {6'h0, gyro1_valid, quat1_valid};
        
        // Sensor 2 Quaternion (MSB,LSB format)
        packet_buffer[16] = quat2_w[15:8];  // W MSB
        packet_buffer[17] = quat2_w[7:0];   // W LSB
        packet_buffer[18] = quat2_x[15:8];  // X MSB
        packet_buffer[19] = quat2_x[7:0];   // X LSB
        packet_buffer[20] = quat2_y[15:8];  // Y MSB
        packet_buffer[21] = quat2_y[7:0];   // Y LSB
        packet_buffer[22] = quat2_z[15:8];  // Z MSB
        packet_buffer[23] = quat2_z[7:0];   // Z LSB
        
        // Sensor 2 Gyroscope (MSB,LSB format)
        packet_buffer[24] = gyro2_x[15:8];  // X MSB
        packet_buffer[25] = gyro2_x[7:0];   // X LSB
        packet_buffer[26] = gyro2_y[15:8];  // Y MSB
        packet_buffer[27] = gyro2_y[7:0];   // Y LSB
        packet_buffer[28] = gyro2_z[15:8];  // Z MSB
        packet_buffer[29] = gyro2_z[7:0];   // Z LSB
        
        // Sensor 2 Flags
        packet_buffer[30] = {6'h0, gyro2_valid, quat2_valid};
        
        // Reserved
        packet_buffer[31] = 8'h00;
    end
    
    // Data ready when either sensor has valid data
    logic data_ready_reg = 1'b0;  // Initialize to 0
    logic has_valid;  // Combinational signal for valid data detection
    logic has_valid_prev = 1'b0;  // Store previous has_valid for edge detection (initialize to 0)
    logic has_valid_prev_reg = 1'b0;  // Register to capture old value before update
    
    assign has_valid = (quat1_valid || gyro1_valid || quat2_valid || gyro2_valid);
    
    always_ff @(posedge clk) begin
        // Update load_prev first (non-blocking, so old value is used in conditions)
        load_prev <= load;
        
        // Check for LOAD edge (acknowledgment) - highest priority
        // load_prev is the OLD value (before the <= assignment above)
        if (load && !load_prev) begin
            // MCU acknowledged - clear data ready
            data_ready_reg <= 1'b0;
            // Set has_valid_prev to current has_valid so we can detect transitions after ack
            has_valid_prev <= has_valid;
            // Update has_valid_prev_reg to track the old value for next cycle
            has_valid_prev_reg <= has_valid_prev;
        end else begin
            // Check conditions using the OLD has_valid_prev value (from has_valid_prev_reg)
            // has_valid_prev_reg contains the value from 2 cycles ago, which is what we need
            // for edge detection (we want to detect when has_valid goes from 0 to 1)
            if (!has_valid) begin
                // No valid data - clear data ready and reset tracking
                data_ready_reg <= 1'b0;
                has_valid_prev <= 1'b0;
                has_valid_prev_reg <= has_valid_prev;  // Update reg to track old value
            end else if (has_valid && !has_valid_prev_reg) begin
                // New data available (valid went from 0 to 1) - set data ready
                // Use has_valid_prev_reg (old value from 2 cycles ago) to detect 0->1 transition
                data_ready_reg <= 1'b1;
                has_valid_prev <= 1'b1;
                has_valid_prev_reg <= has_valid_prev;  // Update reg to track old value
            end else begin
                // Valid data still present (has_valid && has_valid_prev_reg) - keep current state
                // Update has_valid_prev to maintain tracking
                has_valid_prev <= 1'b1;
                has_valid_prev_reg <= has_valid_prev;  // Update reg to track old value
            end
        end
    end
    
    // Done signal: Assert when data is ready
    assign done = data_ready_reg;
    
    // Create a 256-bit shift register from packet buffer (32 bytes * 8 bits)
    logic [255:0] packet_shift_reg;
    
    // SPI transmission: Shift on posedge sck (like aes_spi.sv)
    // Following aes_spi pattern: on first posedge (!wasdone), load AND shift
    // On subsequent posedges (wasdone), shift left
    always_ff @(posedge sck) begin
        if (!wasdone) begin
            // First posedge: load buffer and shift in one operation (like aes_spi)
            // Pack all bytes into shift register: MSB first (packet_buffer[0] is MSB)
            packet_shift_reg <= {
                packet_buffer[0], packet_buffer[1], packet_buffer[2], packet_buffer[3],
                packet_buffer[4], packet_buffer[5], packet_buffer[6], packet_buffer[7],
                packet_buffer[8], packet_buffer[9], packet_buffer[10], packet_buffer[11],
                packet_buffer[12], packet_buffer[13], packet_buffer[14], packet_buffer[15],
                packet_buffer[16], packet_buffer[17], packet_buffer[18], packet_buffer[19],
                packet_buffer[20], packet_buffer[21], packet_buffer[22], packet_buffer[23],
                packet_buffer[24], packet_buffer[25], packet_buffer[26], packet_buffer[27],
                packet_buffer[28], packet_buffer[29], packet_buffer[30], packet_buffer[31],
                sdi  // Shift in SDI on first edge (like aes_spi)
            };
        end else begin
            // Subsequent posedges: shift left (MSB first)
            packet_shift_reg <= {packet_shift_reg[254:0], sdi};
        end
    end
    
    // Track previous done state (for edge detection - like aes_spi)
    // aes_spi uses blocking assignment for immediate update
    always @(negedge sck) begin
        wasdone = done;
        sdodelayed = packet_shift_reg[254];  // Next bit to output (like aes_spi cyphertextcaptured[126])
    end
    
    // SDO output: Following aes_spi pattern exactly
    // When done is first asserted (!wasdone), output MSB before first clock edge
    // After first negedge, wasdone becomes true, so use sdodelayed
    assign sdo = (done & !wasdone) ? packet_buffer[0][7] : sdodelayed;
    
endmodule


